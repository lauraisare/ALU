library verilog;
use verilog.vl_types.all;
entity ALU_test_vlg_vec_tst is
end ALU_test_vlg_vec_tst;
